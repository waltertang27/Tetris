module font_rom ( input [10:0]	addr,
						output [15:0]	data
					 );

	parameter ADDR_WIDTH = 11;
   parameter DATA_WIDTH =  16;
	logic [ADDR_WIDTH-1:0] addr_reg;
				
	// ROM definition				
	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x01 BLOCK TYPE 1
        16'b0011111111111111, // 0   **************
        16'b0011111111111111, // 1   **************
        16'b1100000000000011, // 2 **            **
        16'b1100000000000011, // 3 **            **
        16'b1100000000000011, // 4 **            **
        16'b1100000000000011, // 5 **            **
        16'b1100000000000011, // 6 **            **
        16'b1100000000000011, // 7 **            **
        16'b1100000000000011, // 8 **            **
        16'b1100000000000011, // 9 **            **
        16'b1100000000000011, // a **            **
        16'b1100000000000011, // b **            **
        16'b1100000000000011, // c **            **
        16'b1100000000000011, // d **            **
        16'b1111111111111111, // e ****************
        16'b1111111111111111, // f ****************
         // code x02 BLOCK TYPE 2
        16'b0011111111111111, // 0   **************
        16'b0011111111111111, // 1   **************
        16'b1100001111111111, // 2 **    **********
        16'b1100001111111111, // 3 **    **********
        16'b1100111111111111, // 4 **  ************
        16'b1100111111111111, // 5 **  ************
        16'b1111111111111111, // 6 ****************
        16'b1111111111111111, // 7 ****************
        16'b1111111111111111, // 8 ****************
        16'b1111111111111111, // 9 ****************
        16'b1111111111111111, // a ****************
        16'b1111111111111111, // b ****************
        16'b1111111111111111, // c ****************
        16'b1111111111111111, // d ****************
        16'b1111111111111111, // e ****************
        16'b1111111111111111, // f ****************
         // code x03 TOP LEFT GRID CORNER
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000011111111, // 8         ********
        16'b0000000011111111, // 9         ********
        16'b0000000011111111, // a         ********
        16'b0000000011111111, // b         ********
        16'b0000000011111111, // c         ********
        16'b0000000011111111, // d         ********
        16'b0000000011111111, // e         ********
        16'b0000000011111111, // f         ********
         // code x04 GRID TOP WALL
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b1111111111111111, // 8 ****************
        16'b1111111111111111, // 9 ****************
        16'b1111111111111111, // a ****************
        16'b1111111111111111, // b ****************
        16'b1111111111111111, // c ****************
        16'b1111111111111111, // d ****************
        16'b1111111111111111, // e ****************
        16'b1111111111111111, // f ****************
         // code x05 TOP RIGHT GRID CORNER
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b1111111100000000, // 8 ********
        16'b1111111100000000, // 9 ********
        16'b1111111100000000, // a ********
        16'b1111111100000000, // b ********
        16'b1111111100000000, // c ********
        16'b1111111100000000, // d ********
        16'b1111111100000000, // e ********
        16'b1111111100000000, // f ********
         // code x06 GRID RIGHT WALL
        16'b1111111100000000, // 0 ********
        16'b1111111100000000, // 1 ********
        16'b1111111100000000, // 2 ********
        16'b1111111100000000, // 3 ********
        16'b1111111100000000, // 4 ********
        16'b1111111100000000, // 5 ********
        16'b1111111100000000, // 6 ********
        16'b1111111100000000, // 7 ********
        16'b1111111100000000, // 8 ********
        16'b1111111100000000, // 9 ********
        16'b1111111100000000, // a ********
        16'b1111111100000000, // b ********
        16'b1111111100000000, // c ********
        16'b1111111100000000, // d ********
        16'b1111111100000000, // e ********
        16'b1111111100000000, // f ********
         // code x07 BOTTOM RIGHT GRID CORNER
        16'b1111111100000000, // 0 ********
        16'b1111111100000000, // 1 ********
        16'b1111111100000000, // 2 ********
        16'b1111111100000000, // 3 ********
        16'b1111111100000000, // 4 ********
        16'b1111111100000000, // 5 ********
        16'b1111111100000000, // 6 ********
        16'b1111111100000000, // 7 ********
        16'b0000000000000000, // 8 
        16'b0000000000000000, // 9 
        16'b0000000000000000, // a 
        16'b0000000000000000, // b 
        16'b0000000000000000, // c 
        16'b0000000000000000, // d 
        16'b0000000000000000, // e 
        16'b0000000000000000, // f 
         // code x08 GRID BOTTOM WALL
        16'b1111111111111111, // 0 ****************
        16'b1111111111111111, // 1 ****************
        16'b1111111111111111, // 2 ****************
        16'b1111111111111111, // 3 ****************
        16'b1111111111111111, // 4 ****************
        16'b1111111111111111, // 5 ****************
        16'b1111111111111111, // 6 ****************
        16'b1111111111111111, // 7 ****************
        16'b0000000000000000, // 8 
        16'b0000000000000000, // 9 
        16'b0000000000000000, // a 
        16'b0000000000000000, // b 
        16'b0000000000000000, // c 
        16'b0000000000000000, // d 
        16'b0000000000000000, // e 
        16'b0000000000000000, // f 
         // code x09 BOTTOM LEFT GRID CORNER
        16'b0000000011111111, // 0         ********
        16'b0000000011111111, // 1         ********
        16'b0000000011111111, // 2         ********
        16'b0000000011111111, // 3         ********
        16'b0000000011111111, // 4         ********
        16'b0000000011111111, // 5         ********
        16'b0000000011111111, // 6         ********
        16'b0000000011111111, // 7         ********
        16'b0000000000000000, // 8 
        16'b0000000000000000, // 9 
        16'b0000000000000000, // a 
        16'b0000000000000000, // b 
        16'b0000000000000000, // c 
        16'b0000000000000000, // d 
        16'b0000000000000000, // e 
        16'b0000000000000000, // f 
         // code x0a GRID LEFT WALL
        16'b0000000011111111, // 0         ********
        16'b0000000011111111, // 1         ********
        16'b0000000011111111, // 2         ********
        16'b0000000011111111, // 3         ********
        16'b0000000011111111, // 4         ********
        16'b0000000011111111, // 5         ********
        16'b0000000011111111, // 6         ********
        16'b0000000011111111, // 7         ********
        16'b0000000011111111, // 8         ********
        16'b0000000011111111, // 9         ********
        16'b0000000011111111, // a         ********
        16'b0000000011111111, // b         ********
        16'b0000000011111111, // c         ********
        16'b0000000011111111, // d         ********
        16'b0000000011111111, // e         ********
        16'b0000000011111111, // f         ********
         // code x0b SMALL TOP LEFT CORNER
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000011, // e               **
        16'b0000000000000011, // f               **
         // code x0c SMALL TOP WALL
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b1111111111111111, // e ****************
        16'b1111111111111111, // f ****************
         // code x0d SMALL TOP RIGHT CORNER
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b1100000000000000, // e **
        16'b1100000000000000, // f **
         // code x0e SMALL RIGHT WALL
        16'b1100000000000000, // 0 **
        16'b1100000000000000, // 1 **
        16'b1100000000000000, // 2 **
        16'b1100000000000000, // 3 **
        16'b1100000000000000, // 4 **
        16'b1100000000000000, // 5 **
        16'b1100000000000000, // 6 **
        16'b1100000000000000, // 7 **
        16'b1100000000000000, // 8 **
        16'b1100000000000000, // 9 **
        16'b1100000000000000, // a **
        16'b1100000000000000, // b **
        16'b1100000000000000, // c **
        16'b1100000000000000, // d **
        16'b1100000000000000, // e **
        16'b1100000000000000, // f **
         // code x0f SMALL BOTTOM RIGHT CORNER
        16'b1100000000000000, // 0 **
        16'b1100000000000000, // 1 **
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x10 SMALL BOTTOM WALL
        16'b1111111111111111, // 0 ****************
        16'b1111111111111111, // 1 ****************
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x11 SMALL BOTTOM LEFT CORNER
        16'b0000000000000011, // 0               **
        16'b0000000000000011, // 1               **
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x12 SMALL LEFT WALL
        16'b0000000000000011, // 0               **
        16'b0000000000000011, // 1               **
        16'b0000000000000011, // 2               **
        16'b0000000000000011, // 3               **
        16'b0000000000000011, // 4               **
        16'b0000000000000011, // 5               **
        16'b0000000000000011, // 6               **
        16'b0000000000000011, // 7               **
        16'b0000000000000011, // 8               **
        16'b0000000000000011, // 9               **
        16'b0000000000000011, // a               **
        16'b0000000000000011, // b               **
        16'b0000000000000011, // c               **
        16'b0000000000000011, // d               **
        16'b0000000000000011, // e               **
        16'b0000000000000011, // f               **
         // code x13
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x14
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x15
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x16
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x17
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x18
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x19
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x1a
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x1b
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x1c
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x1d
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x1e
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x1f
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x20
        16'b0000000000000000, // 0
        16'b0111111111111110, // 1 **************
        16'b0111111111111110, // 2 **************
        16'b0111111111111110, // 3 **************
        16'b0111100000011110, // 4 ****      ****
        16'b0111100000011110, // 5 ****      ****
        16'b0111100000011110, // 6 ****      ****
        16'b0111111111111110, // 7 **************
        16'b0111111111111110, // 8 **************
        16'b0111111111111110, // 9 **************
        16'b0111100000011110, // a ****      ****
        16'b0111100000011110, // b ****      ****
        16'b0111100000011110, // c ****      ****
        16'b0111100000011110, // d ****      ****
        16'b0111100000011110, // e ****      ****
        16'b0000000000000000, // f
         // code x21
        16'b0000000000000000, // 0
        16'b0111111111111100, // 1 *************
        16'b0111111111111110, // 2 **************
        16'b0111111111111110, // 3 **************
        16'b0111100000011110, // 4 ****      ****
        16'b0111100000011110, // 5 ****      ****
        16'b0111111111111110, // 6 **************
        16'b0111111111111110, // 7 **************
        16'b0111111111111100, // 8 *************
        16'b0111100000011100, // 9 ****      ***
        16'b0111100000011110, // a ****      ****
        16'b0111100000011110, // b ****      ****
        16'b0111111111111110, // c **************
        16'b0111111111111110, // d **************
        16'b0111111111111100, // e *************
        16'b0000000000000000, // f
         // code x22
        16'b0000000000000000, // 0
        16'b0111111111111110, // 1 **************
        16'b0111111111111110, // 2 **************
        16'b0111111111111110, // 3 **************
        16'b0111100000000000, // 4 ****
        16'b0111100000000000, // 5 ****
        16'b0111100000000000, // 6 ****
        16'b0111100000000000, // 7 ****
        16'b0111100000000000, // 8 ****
        16'b0111100000000000, // 9 ****
        16'b0111100000000000, // a ****
        16'b0111100000000000, // b ****
        16'b0111111111111110, // c **************
        16'b0111111111111110, // d **************
        16'b0111111111111110, // e **************
        16'b0000000000000000, // f
         // code x23
        16'b0000000000000000, // 0
        16'b0111111111111100, // 1 *************
        16'b0111111111111110, // 2 **************
        16'b0111111111111110, // 3 **************
        16'b0111100000011110, // 4 ****      ****
        16'b0111100000011110, // 5 ****      ****
        16'b0111100000011110, // 6 ****      ****
        16'b0111100000011110, // 7 ****      ****
        16'b0111100000011110, // 8 ****      ****
        16'b0111100000011110, // 9 ****      ****
        16'b0111100000011110, // a ****      ****
        16'b0111100000011110, // b ****      ****
        16'b0111111111111110, // c **************
        16'b0111111111111110, // d **************
        16'b0111111111111100, // e *************
        16'b0000000000000000, // f
         // code x24
        16'b0000000000000000, // 0
        16'b0111111111111110, // 1 **************
        16'b0111111111111110, // 2 **************
        16'b0111111111111110, // 3 **************
        16'b0111100000000000, // 4 ****
        16'b0111100000000000, // 5 ****
        16'b0111111111111100, // 6 *************
        16'b0111111111111100, // 7 *************
        16'b0111111111111100, // 8 *************
        16'b0111100000000000, // 9 ****
        16'b0111100000000000, // a ****
        16'b0111100000000000, // b ****
        16'b0111111111111110, // c **************
        16'b0111111111111110, // d **************
        16'b0111111111111110, // e **************
        16'b0000000000000000, // f
         // code x25
        16'b0000000000000000, // 0
        16'b0111111111111110, // 1 **************
        16'b0111111111111110, // 2 **************
        16'b0111111111111110, // 3 **************
        16'b0111100000000000, // 4 ****
        16'b0111100000000000, // 5 ****
        16'b0111111111111100, // 6 *************
        16'b0111111111111100, // 7 *************
        16'b0111111111111100, // 8 *************
        16'b0111100000000000, // 9 ****
        16'b0111100000000000, // a ****
        16'b0111100000000000, // b ****
        16'b0111100000000000, // c ****
        16'b0111100000000000, // d ****
        16'b0111100000000000, // e ****
        16'b0000000000000000, // f
         // code x26
        16'b0000000000000000, // 0
        16'b0111111111111110, // 1 **************
        16'b0111111111111110, // 2 **************
        16'b0111111111111110, // 3 **************
        16'b0111100000000000, // 4 ****
        16'b0111100000000000, // 5 ****
        16'b0111100000000000, // 6 ****
        16'b0111100000000000, // 7 ****
        16'b0111100001111110, // 8 ****    ******
        16'b0111100001111110, // 9 ****    ******
        16'b0111100000011110, // a ****      ****
        16'b0111100000011110, // b ****      ****
        16'b0111111111111110, // c **************
        16'b0111111111111110, // d **************
        16'b0111111111111110, // e **************
        16'b0000000000000000, // f
         // code x27
        16'b0000000000000000, // 0
        16'b0111100000011110, // 1 ****      ****
        16'b0111100000011110, // 2 ****      ****
        16'b0111100000011110, // 3 ****      ****
        16'b0111100000011110, // 4 ****      ****
        16'b0111100000011110, // 5 ****      ****
        16'b0111111111111110, // 6 **************
        16'b0111111111111110, // 7 **************
        16'b0111111111111110, // 8 **************
        16'b0111111111111110, // 9 **************
        16'b0111100000011110, // a ****      ****
        16'b0111100000011110, // b ****      ****
        16'b0111100000011110, // c ****      ****
        16'b0111100000011110, // d ****      ****
        16'b0111100000011110, // e ****      ****
        16'b0000000000000000, // f
         // code x28
        16'b0000000000000000, // 0
        16'b0111111111111110, // 1 **************
        16'b0111111111111110, // 2 **************
        16'b0111111111111110, // 3 **************
        16'b0000001111000000, // 4      ****
        16'b0000001111000000, // 5      ****
        16'b0000001111000000, // 6      ****
        16'b0000001111000000, // 7      ****
        16'b0000001111000000, // 8      ****
        16'b0000001111000000, // 9      ****
        16'b0000001111000000, // a      ****
        16'b0000001111000000, // b      ****
        16'b0111111111111110, // c **************
        16'b0111111111111110, // d **************
        16'b0111111111111110, // e **************
        16'b0000000000000000, // f
         // code x29
        16'b0000000000000000, // 0
        16'b0111111111111110, // 1 **************
        16'b0111111111111110, // 2 **************
        16'b0111111111111110, // 3 **************
        16'b0000000011110000, // 4        ****
        16'b0000000011110000, // 5        ****
        16'b0000000011110000, // 6        ****
        16'b0000000011110000, // 7        ****
        16'b0000000011110000, // 8        ****
        16'b0000000011110000, // 9        ****
        16'b0111000011110000, // a ***    ****
        16'b0111000011110000, // b ***    ****
        16'b0111111111110000, // c ***********
        16'b0111111111110000, // d ***********
        16'b0111111111110000, // e ***********
        16'b0000000000000000, // f
         // code x2a
        16'b0000000000000000, // 0
        16'b0111100000001110, // 1 ****       ***
        16'b0111100000001110, // 2 ****       ***
        16'b0111100000111000, // 3 ****     ***
        16'b0111100000111000, // 4 ****     ***
        16'b0111100111100000, // 5 ****  ****
        16'b0111100111100000, // 6 ****  ****
        16'b0111111110000000, // 7 ********
        16'b0111111110000000, // 8 ********
        16'b0111100111100000, // 9 ****  ****
        16'b0111100111100000, // a ****  ****
        16'b0111100001111000, // b ****    ****
        16'b0111100001111000, // c ****    ****
        16'b0111100000011110, // d ****      ****
        16'b0111100000011110, // e ****      ****
        16'b0000000000000000, // f
         // code x2b
        16'b0000000000000000, // 0
        16'b0111100000000000, // 1 ****
        16'b0111100000000000, // 2 ****
        16'b0111100000000000, // 3 ****
        16'b0111100000000000, // 4 ****
        16'b0111100000000000, // 5 ****
        16'b0111100000000000, // 6 ****
        16'b0111100000000000, // 7 ****
        16'b0111100000000000, // 8 ****
        16'b0111100000000000, // 9 ****
        16'b0111100000000000, // a ****
        16'b0111100000000000, // b ****
        16'b0111111111111110, // c **************
        16'b0111111111111110, // d **************
        16'b0111111111111110, // e **************
        16'b0000000000000000, // f
         // code x2c
        16'b0000000000000000, // 0
        16'b0111100000011110, // 1 ****      ****
        16'b0111100000011110, // 2 ****      ****
        16'b0111100000011110, // 3 ****      ****
        16'b0111111001111110, // 4 ******  ******
        16'b0111111001111110, // 5 ******  ******
        16'b0111111111111110, // 6 **************
        16'b0111111111111110, // 7 **************
        16'b0111100110011110, // 8 ****  **  ****
        16'b0111100110011110, // 9 ****  **  ****
        16'b0111100000011110, // a ****      ****
        16'b0111100000011110, // b ****      ****
        16'b0111100000011110, // c ****      ****
        16'b0111100000011110, // d ****      ****
        16'b0111100000011110, // e ****      ****
        16'b0000000000000000, // f
         // code x2d
        16'b0000000000000000, // 0
        16'b0111100000011110, // 1 ****      ****
        16'b0111100000011110, // 2 ****      ****
        16'b0111100000011110, // 3 ****      ****
        16'b0111111000011110, // 4 ******    ****
        16'b0111111000011110, // 5 ******    ****
        16'b0111111110011110, // 6 ********  ****
        16'b0111111110011110, // 7 ********  ****
        16'b0111100111111110, // 8 ****  ********
        16'b0111100111111110, // 9 ****  ********
        16'b0111100001111110, // a ****    ******
        16'b0111100001111110, // b ****    ******
        16'b0111100000011110, // c ****      ****
        16'b0111100000011110, // d ****      ****
        16'b0111100000011110, // e ****      ****
        16'b0000000000000000, // f
         // code x2e
        16'b0000000000000000, // 0
        16'b0111111111111110, // 1 **************
        16'b0111111111111110, // 2 **************
        16'b0111111111111110, // 3 **************
        16'b0111100000011110, // 4 ****      ****
        16'b0111100000011110, // 5 ****      ****
        16'b0111100000011110, // 6 ****      ****
        16'b0111100000011110, // 7 ****      ****
        16'b0111100000011110, // 8 ****      ****
        16'b0111100000011110, // 9 ****      ****
        16'b0111100000011110, // a ****      ****
        16'b0111100000011110, // b ****      ****
        16'b0111111111111110, // c **************
        16'b0111111111111110, // d **************
        16'b0111111111111110, // e **************
        16'b0000000000000000, // f
         // code x2f
        16'b0000000000000000, // 0
        16'b0111111111111000, // 1 ************
        16'b0111111111111110, // 2 **************
        16'b0111111111111110, // 3 **************
        16'b0111100000011110, // 4 ****      ****
        16'b0111100000011110, // 5 ****      ****
        16'b0111111111111110, // 6 **************
        16'b0111111111111000, // 7 ************
        16'b0111111111111000, // 8 ************
        16'b0111100000000000, // 9 ****
        16'b0111100000000000, // a ****
        16'b0111100000000000, // b ****
        16'b0111100000000000, // c ****
        16'b0111100000000000, // d ****
        16'b0111100000000000, // e ****
        16'b0000000000000000, // f
         // code x30
        16'b0000000000000000, // 0
        16'b0111111111111110, // 1 **************
        16'b0111111111111110, // 2 **************
        16'b0111111111111110, // 3 **************
        16'b0111000000000110, // 4 ***         **
        16'b0111000000000110, // 5 ***         **
        16'b0111000000000110, // 6 ***         **
        16'b0111000000000110, // 7 ***         **
        16'b0111000000000110, // 8 ***         **
        16'b0111000000000110, // 9 ***         **
        16'b0111000011000110, // a ***    **   **
        16'b0111000011000110, // b ***    **   **
        16'b0111111111111000, // c ************
        16'b0111111111111000, // d ************
        16'b0000000000011110, // e           ****
        16'b0000000000000000, // f
         // code x31
        16'b0000000000000000, // 0
        16'b0111111111111000, // 1 ************
        16'b0111111111111110, // 2 **************
        16'b0111111111111110, // 3 **************
        16'b0111100000011110, // 4 ****      ****
        16'b0111100000011110, // 5 ****      ****
        16'b0111111111111110, // 6 **************
        16'b0111111111111000, // 7 ************
        16'b0111111111111000, // 8 ************
        16'b0111100000011110, // 9 ****      ****
        16'b0111100000011110, // a ****      ****
        16'b0111100000011110, // b ****      ****
        16'b0111100000011110, // c ****      ****
        16'b0111100000011110, // d ****      ****
        16'b0111100000011110, // e ****      ****
        16'b0000000000000000, // f
         // code x32
        16'b0000000000000000, // 0
        16'b0111111111111110, // 1 **************
        16'b0111111111111110, // 2 **************
        16'b0111111111111110, // 3 **************
        16'b0111100000000000, // 4 ****
        16'b0111100000000000, // 5 ****
        16'b0111111111111110, // 6 **************
        16'b0111111111111110, // 7 **************
        16'b0111111111111110, // 8 **************
        16'b0000000000011110, // 9           ****
        16'b0000000000011110, // a           ****
        16'b0000000000011110, // b           ****
        16'b0111111111111110, // c **************
        16'b0111111111111110, // d **************
        16'b0111111111111110, // e **************
        16'b0000000000000000, // f
         // code x33
        16'b0000000000000000, // 0
        16'b0111111111111110, // 1 **************
        16'b0111111111111110, // 2 **************
        16'b0111111111111110, // 3 **************
        16'b0000001111000000, // 4      ****
        16'b0000001111000000, // 5      ****
        16'b0000001111000000, // 6      ****
        16'b0000001111000000, // 7      ****
        16'b0000001111000000, // 8      ****
        16'b0000001111000000, // 9      ****
        16'b0000001111000000, // a      ****
        16'b0000001111000000, // b      ****
        16'b0000001111000000, // c      ****
        16'b0000001111000000, // d      ****
        16'b0000001111000000, // e      ****
        16'b0000000000000000, // f
         // code x34
        16'b0000000000000000, // 0
        16'b0111100000011110, // 1 ****      ****
        16'b0111100000011110, // 2 ****      ****
        16'b0111100000011110, // 3 ****      ****
        16'b0111100000011110, // 4 ****      ****
        16'b0111100000011110, // 5 ****      ****
        16'b0111100000011110, // 6 ****      ****
        16'b0111100000011110, // 7 ****      ****
        16'b0111100000011110, // 8 ****      ****
        16'b0111100000011110, // 9 ****      ****
        16'b0111100000011110, // a ****      ****
        16'b0111100000011110, // b ****      ****
        16'b0111111111111110, // c **************
        16'b0111111111111110, // d **************
        16'b0111111111111110, // e **************
        16'b0000000000000000, // f
         // code x35
        16'b0000000000000000, // 0
        16'b0111100000011110, // 1 ****      ****
        16'b0111100000011110, // 2 ****      ****
        16'b0111100000011110, // 3 ****      ****
        16'b0111100000011110, // 4 ****      ****
        16'b0111100000011110, // 5 ****      ****
        16'b0111100000011110, // 6 ****      ****
        16'b0111100000011110, // 7 ****      ****
        16'b0001111001111000, // 8   ****  ****
        16'b0001111001111000, // 9   ****  ****
        16'b0001111001111000, // a   ****  ****
        16'b0001111001111000, // b   ****  ****
        16'b0000011111100000, // c     ******
        16'b0000011111100000, // d     ******
        16'b0000011111100000, // e     ******
        16'b0000000000000000, // f
         // code x36
        16'b0000000000000000, // 0
        16'b0111100000011110, // 1 ****      ****
        16'b0111100000011110, // 2 ****      ****
        16'b0111100000011110, // 3 ****      ****
        16'b0111100000011110, // 4 ****      ****
        16'b0111100000011110, // 5 ****      ****
        16'b0111100000011110, // 6 ****      ****
        16'b0111100110011110, // 7 ****  **  ****
        16'b0111100110011110, // 8 ****  **  ****
        16'b0111111111111110, // 9 **************
        16'b0111111111111110, // a **************
        16'b0111111001111110, // b ******  ******
        16'b0111111001111110, // c ******  ******
        16'b0111100000011110, // d ****      ****
        16'b0111100000011110, // e ****      ****
        16'b0000000000000000, // f
         // code x37
        16'b0000000000000000, // 0 
        16'b0111100000011110, // 1 ****      ****
        16'b0111100000011110, // 2 ****      ****
        16'b0111100000011110, // 3 ****      ****
        16'b0001111001111000, // 4   ****  ****
        16'b0001111001111000, // 5   ****  ****
        16'b0000011111100000, // 6     ******
        16'b0000011111100000, // 7     ******
        16'b0000011111100000, // 8     ******
        16'b0000011111100000, // 9     ******
        16'b0001111001111000, // a   ****  ****
        16'b0001111001111000, // b   ****  ****
        16'b0111100000011110, // c ****      ****
        16'b0111100000011110, // d ****      ****
        16'b0111100000011110, // e ****      ****
        16'b0000000000000000, // f
         // code x38
        16'b0000000000000000, // 0
        16'b0111100000011110, // 1 ****      ****
        16'b0111100000011110, // 2 ****      ****
        16'b0111100000011110, // 3 ****      ****
        16'b0111100000011110, // 4 ****      ****
        16'b0111111001111110, // 5 ******  ******
        16'b0111111001111110, // 6 ******  ******
        16'b0001111111111000, // 7   **********
        16'b0001111111111000, // 8   **********
        16'b0000011111100000, // 9     ******
        16'b0000011111100000, // a     ******
        16'b0000011111100000, // b     ******
        16'b0000011111100000, // c     ******
        16'b0000011111100000, // d     ******
        16'b0000011111100000, // e     ******
        16'b0000000000000000, // f
         // code x39
        16'b0000000000000000, // 0
        16'b0111111111111110, // 1 **************
        16'b0111111111111110, // 2 **************
        16'b0111111111111110, // 3 **************
        16'b0000000001111000, // 4         ****
        16'b0000000001111000, // 5         ****
        16'b0000000111100000, // 6       ****
        16'b0000000111100000, // 7       ****
        16'b0000011110000000, // 8     ****
        16'b0000011110000000, // 9     ****
        16'b0001111000000000, // a   ****
        16'b0001111000000000, // b   ****
        16'b0111111111111110, // c **************
        16'b0111111111111110, // d **************
        16'b0111111111111110, // e **************
        16'b0000000000000000, // f
         // code x3a
        16'b0000000000000000, // 0
        16'b0000001111000000, // 1      ****
        16'b0000001111000000, // 2      ****
        16'b0000001111000000, // 3      ****
        16'b0000001111000000, // 4      ****
        16'b0000001111000000, // 5      ****
        16'b0000001111000000, // 6      ****
        16'b0000001111000000, // 7      ****
        16'b0000001111000000, // 8      ****
        16'b0000001111000000, // 9      ****
        16'b0000001111000000, // a      ****
        16'b0000001111000000, // b      ****
        16'b0000001111000000, // c      ****
        16'b0000001111000000, // d      ****
        16'b0000001111000000, // e      ****
        16'b0000000000000000, // f
         // code x3b
        16'b0000000000000000, // 0
        16'b0111111111111110, // 1 **************
        16'b0111111111111110, // 2 **************
        16'b0111111111111110, // 3 **************
        16'b0000000000011110, // 4           ****
        16'b0000000000011110, // 5           ****
        16'b0111111111111110, // 6 **************
        16'b0111111111111110, // 7 **************
        16'b0111111111111110, // 8 **************
        16'b0111100000000000, // 9 ****
        16'b0111100000000000, // a ****
        16'b0111100000000000, // b ****
        16'b0111111111111110, // c **************
        16'b0111111111111110, // d **************
        16'b0111111111111110, // e **************
        16'b0000000000000000, // f
         // code x3c
        16'b0000000000000000, // 0
        16'b0111111111111110, // 1 **************
        16'b0111111111111110, // 2 **************
        16'b0111111111111110, // 3 **************
        16'b0000000000011110, // 4           ****
        16'b0000000000011110, // 5           ****
        16'b0111111111111110, // 6 **************
        16'b0111111111111110, // 7 **************
        16'b0111111111111110, // 8 **************
        16'b0000000000011110, // 9           ****
        16'b0000000000011110, // a           ****
        16'b0000000000011110, // b           ****
        16'b0111111111111110, // c **************
        16'b0111111111111110, // d **************
        16'b0111111111111110, // e **************
        16'b0000000000000000, // f
         // code x3d
        16'b0000000000000000, // 0
        16'b0111100000011110, // 1 ****      ****
        16'b0111100000011110, // 2 ****      ****
        16'b0111100000011110, // 3 ****      ****
        16'b0111100000011110, // 4 ****      ****
        16'b0111100000011110, // 5 ****      ****
        16'b0111111111111110, // 6 **************
        16'b0111111111111110, // 7 **************
        16'b0111111111111110, // 8 **************
        16'b0111111111111110, // 9 **************
        16'b0000000000011110, // a           ****
        16'b0000000000011110, // b           ****
        16'b0000000000011110, // c           ****
        16'b0000000000011110, // d           ****
        16'b0000000000011110, // e           ****
        16'b0000000000000000, // f
         // code x3e
        16'b0000000000000000, // 0
        16'b0111111111111110, // 1 **************
        16'b0111111111111110, // 2 **************
        16'b0111111111111110, // 3 **************
        16'b0111100000000000, // 4 ****
        16'b0111100000000000, // 5 ****
        16'b0111111111111110, // 6 **************
        16'b0111111111111110, // 7 **************
        16'b0111111111111110, // 8 **************
        16'b0000000000011110, // 9           ****
        16'b0000000000011110, // a           ****
        16'b0000000000011110, // b           ****
        16'b0111111111111110, // c **************
        16'b0111111111111110, // d **************
        16'b0111111111111110, // e **************
        16'b0000000000000000, // f
         // code x3f
        16'b0000000000000000, // 0
        16'b0111111111111110, // 1 **************
        16'b0111111111111110, // 2 **************
        16'b0111111111111110, // 3 **************
        16'b0111100000000000, // 4 ****
        16'b0111100000000000, // 5 ****
        16'b0111111111111110, // 6 **************
        16'b0111111111111110, // 7 **************
        16'b0111111111111110, // 8 **************
        16'b0111100000011110, // 9 ****      ****
        16'b0111100000011110, // a ****      ****
        16'b0111100000011110, // b ****      ****
        16'b0111111111111110, // c **************
        16'b0111111111111110, // d **************
        16'b0111111111111110, // e **************
        16'b0000000000000000, // f
         // code x40
        16'b0000000000000000, // 0
        16'b0111111111111110, // 1 **************
        16'b0111111111111110, // 2 **************
        16'b0111111111111110, // 3 **************
        16'b0000000000011110, // 4           ****
        16'b0000000000011110, // 5           ****
        16'b0000000000011110, // 6           ****
        16'b0000000000011110, // 7           ****
        16'b0000000000011110, // 8           ****
        16'b0000000000011110, // 9           ****
        16'b0000000000011110, // a           ****
        16'b0000000000011110, // b           ****
        16'b0000000000011110, // c           ****
        16'b0000000000011110, // d           ****
        16'b0000000000011110, // e           ****
        16'b0000000000000000, // f
         // code x41
        16'b0000000000000000, // 0
        16'b0111111111111110, // 1 **************
        16'b0111111111111110, // 2 **************
        16'b0111111111111110, // 3 **************
        16'b0111100000011110, // 4 ****      ****
        16'b0111100000011110, // 5 ****      ****
        16'b0111111111111110, // 6 **************
        16'b0111111111111110, // 7 **************
        16'b0111111111111110, // 8 **************
        16'b0111100000011110, // 9 ****      ****
        16'b0111100000011110, // a ****      ****
        16'b0111100000011110, // b ****      ****
        16'b0111111111111110, // c **************
        16'b0111111111111110, // d **************
        16'b0111111111111110, // e **************
        16'b0000000000000000, // f
         // code x42
        16'b0000000000000000, // 0
        16'b0111111111111110, // 1 **************
        16'b0111111111111110, // 2 **************
        16'b0111111111111110, // 3 **************
        16'b0111100000011110, // 4 ****      ****
        16'b0111100000011110, // 5 ****      ****
        16'b0111111111111110, // 6 **************
        16'b0111111111111110, // 7 **************
        16'b0111111111111110, // 8 **************
        16'b0000000000011110, // 9           ****
        16'b0000000000011110, // a           ****
        16'b0000000000011110, // b           ****
        16'b0000000000011110, // c           ****
        16'b0000000000011110, // d           ****
        16'b0000000000011110, // e           ****
        16'b0000000000000000, // f
         // code x43
        16'b0000000000000000, // 0
        16'b0111111111111110, // 1 **************
        16'b0111111111111110, // 2 **************
        16'b0111111111111110, // 3 **************
        16'b0111100000011110, // 4 ****      ****
        16'b0111100000011110, // 5 ****      ****
        16'b0111100110011110, // 6 ****  **  ****
        16'b0111100110011110, // 7 ****  **  ****
        16'b0111100110011110, // 8 ****  **  ****
        16'b0111100110011110, // 9 ****  **  ****
        16'b0111100000011110, // a ****      ****
        16'b0111100000011110, // b ****      ****
        16'b0111111111111110, // c **************
        16'b0111111111111110, // d **************
        16'b0111111111111110, // e **************
        16'b0000000000000000, // f
         // code x44
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0011110000000000, // 2  ****
        16'b0011110000000000, // 3  ****
        16'b0011110000000000, // 4  ****
        16'b0011110000000000, // 5  ****
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0011110000000000, // a  ****
        16'b0011110000000000, // b  ****
        16'b0011110000000000, // c  ****
        16'b0011110000000000, // d  ****
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x45
        16'b0000000000000000, // 0
        16'b0011110000000000, // 1  ****
        16'b0011110000000000, // 2  ****
        16'b0011110000000000, // 3  ****
        16'b0011110000000000, // 4  ****
        16'b0011110000000000, // 5  ****
        16'b0011110000000000, // 6  ****
        16'b0011110000000000, // 7  ****
        16'b0011110000000000, // 8  ****
        16'b0011110000000000, // 9  ****
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0011110000000000, // c  ****
        16'b0011110000000000, // d  ****
        16'b0011110000000000, // e  ****
        16'b0000000000000000, // f
         // code x46
        16'b0000000000000000, // 0
        16'b0111111111111110, // 1 **************
        16'b0111111111111110, // 2 **************
        16'b0111111111111110, // 3 **************
        16'b0111100000011110, // 4 ****      ****
        16'b0111100000011110, // 5 ****      ****
        16'b0111100111111110, // 6 ****  ********
        16'b0111100111111110, // 7 ****  ********
        16'b0000000111100000, // 8       ****
        16'b0000000111100000, // 9       ****
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000111100000, // c       ****
        16'b0000000111100000, // d       ****
        16'b0000000111100000, // e       ****
        16'b0000000000000000, // f
         // code x47
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x48
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x49
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x4a
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x4b
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x4c
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x4d
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x4e
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x4f
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x50
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x510
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x52
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x53
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x54
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x55
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x56
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x57
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
        
         // code x58
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x59
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x5a
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x5b
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x5c
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x5d
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x5e
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x5f
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x60
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x61
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x62
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x63
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x64
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x65
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x66
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x67
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x68
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x69
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x6a
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x6b
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x6c
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x6d
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x6e
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x6f
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x70
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x71
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x72
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x73
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x74
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x75
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x76
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x77
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x78
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x79
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x7a
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x7b
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x7c
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x7d
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x7e
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
         // code x7f
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 3
        16'b0000000000000000, // 4
        16'b0000000000000000, // 5
        16'b0000000000000000, // 6
        16'b0000000000000000, // 7
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000, // f
        };

	assign data = ROM[addr];

endmodule  